module sysdeps

pub fn example() {
	return
}
