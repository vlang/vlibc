module main

#flag -ffreestanding
#flag -c

fn main() {
	return
}
