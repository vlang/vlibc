module main

import sysdeps

#flag -ffreestanding
#flag -c

fn main() {
	sysdeps.example()
}
